
module count4 (
    input clock,
    # signals
    input enable,
    input reset,
    output wire [3:0] count
)