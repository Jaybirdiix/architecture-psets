
module count4 (
    input clock,
    # signal
    input enable,
)