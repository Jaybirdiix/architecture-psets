
module count4 (
    input clock,
    
)