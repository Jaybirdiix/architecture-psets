
module count4 (
    input clock,
    input enable,
)