
module count4 (
    input clock,
    # signals
    input enable,
)