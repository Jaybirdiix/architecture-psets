
module count4 (
    input clock,
    // signals
    input enable,
    input reset,
    // output
    output wire [3:0] count
)

reg [3:0]

endmodule